//-------------------------------------------------------------
//  Tech Task 1 - Xilinx
//  Clock Period Package
//  Author : Sheshu Ramanandan : krsheshu@gmail.com
//-------------------------------------------------------------

package clock_period_pkg;

    parameter CLKPERIOD_NS = 8.196       ;   // 122MHz

endpackage
